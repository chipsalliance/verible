module instance_parameters;
  bar #(4, 8) baz;
endmodule
