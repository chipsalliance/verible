module truncated_numeric_literal;
  assign a = 4'h1F;
endmodule
