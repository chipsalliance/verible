// Copyright 2020 Google LLC.
// SPDX-License-Identifier: Apache-2.0

//- @bad_goal ref _
module bad_goal;
endmodule
