class my_class3;
    static int x;

    static function int my_fun();
        return x;
    endfunction
endclass
