module 654foo;  // lexer should reject invalid identifier
endmodule
