// 'localparams' should only be declared within modules' and classes' definition bodies.
localparam int Foo = 1;
