// Macro name must be styled with all capital letters, underscores, or digits.
`define Foo
