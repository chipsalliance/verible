//- @MyClassIncludedFile1 defines/binding MyClassIncludedFile1
class MyClassIncludedFile1;
    //- @var6 defines/binding Var6
    static int var6;

    //- @my_fun1 defines/binding MyFun1
    static function int my_fun1();
        return 1;
    endfunction
endclass