// Copyright 2020 Google LLC.
// SPDX-License-Identifier: Apache-2.0

//- @"\"D.svh\"" ref/includes Dsvh
//- Dsvh.node/kind file
`include "D.svh"

//- @E defines/binding _
//- @D ref D
localparam E = D;
