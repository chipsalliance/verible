module forbid_negative_array_dim ();
  reg [-1 : 0] x;
endmodule
