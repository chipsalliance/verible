module forbid_consecutive_null_statements;
    ;; // [Style: consecutive-null-statements] [forbid-consecutive-null-statements]
endmodule
