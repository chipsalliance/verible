// Expects all function parameters to explicitly define a storage type.
function automatic int foo(bar = 1);
endfunction
