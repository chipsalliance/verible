// Expect the parameter to explicitly define a storage type
parameter Bar = 1;
