//- @B defines/binding B
//- @A ref A
localparam B = A + 1;
