module instance_ports;
  bar baz(x, y);
endmodule
