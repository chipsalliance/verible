module generate_label_module;
  generate if (foo) begin
    baz bam;
  end
  endgenerate
endmodule
