// All unions should be typedef'd
union {
    bit [8:0] flags;
    int val;
} custom;
