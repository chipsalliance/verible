// Each file should have only one module

module one_module_per_file;
// module name must be the same as file name
endmodule
module second;
endmodule
