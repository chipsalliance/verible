// Expand blocks with two or more expressions
//
// gh_issue: https://github.com/google/verible/issues/445

constraint param_c {a_param == 0; d_param == 0;}
