// Struct names should be lower_snake_case and end with '_t'
typedef struct packed{
    int x, y;
} camelStruct;
