module explicit_begin ();
    always_comb
        a = 1;
endmodule
