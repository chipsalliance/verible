// This case statement is missing a default case
function automatic int foo (input bit in);
  case (in)
    1: return 0;
  endcase
endfunction
