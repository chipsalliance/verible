// Missing explicit lifetime declaration
task foo();
endtask
