// Copyright 2020 Google LLC.
// SPDX-License-Identifier: Apache-2.0

//- @A defines/binding A
localparam A = 1;
