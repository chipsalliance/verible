// verilog_syntax: parse-as-module-body
// verilog_lint: waive legacy-generate-region
generate if (foo) begin
  baz bam;
end
endgenerate
