// All structs should be typedef'd
struct {
    int x,y;
} point;
