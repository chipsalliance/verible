// Interface names should be lower_snake_case and end with _if
interface fooBar;
endinterface
