// 'parameters' should only be declared within packages or parameterized modules/classes.
module proper_parameter_declaration;
  parameter int Bar = 1;
endmodule
