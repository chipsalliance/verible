// All enum declarations should be named with typedef
enum logic [1:0] {
    IsIdle,
    IsRunning,
    IsBlocked
} a_status;
