package endif_comment;
`ifdef FOOBAR
  parameter int P = 4;
`endif
endpackage
