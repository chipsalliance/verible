// Copyright 2020 Google LLC.
// SPDX-License-Identifier: Apache-2.0

//- @D defines/binding D
localparam D = 1;
