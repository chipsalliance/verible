module undersized_binary_literal;
  localparam logic [1:0] Foo = 2'b1;
endmodule
