module foo;
endmodule
