module	tabs; // tabs bad!
endmodule
