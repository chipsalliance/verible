class foo;
  function void bar();
    void'(randomize());
  endfunction
endclass
