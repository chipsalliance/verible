module forbid_implicit_declarations;
  assign a1 = 1'b0; // [Style: implicit-declarations] [forbid-implicit-declarations]
endmodule
