module wrong_module_name;
endmodule
