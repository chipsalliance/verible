// Expects all task parameters to explicitly define a storage type.
task automatic foo(bar = 1);
endtask
