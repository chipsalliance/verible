class foo;
  task bar;
    `uvm_warning("use uvm_error or uvm_info")
  endtask
endclass
