// Expects module port 'helloWorld' to follow lower_snake_case naming convention.
module signal_name_style(input bit helloWorld);
endmodule
