module generate_label_prefix;
  genvar i;
  for (i = 0; i < 5; ++i) begin : invalid_label
  end
endmodule
