// Interface names should be lower_snake_case and end with _if
typedef virtual interface foo barBaz;
