//- @A defines/binding A
localparam A = 1;
