// Expected parameter name, "Hello_World" to follow UpperCamelCase or ALL_CAPS naming convention.
parameter int Hello_World = 1;
