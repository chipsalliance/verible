// Expected localparam name, "Hello_World" to follow UpperCamelCase
// naming convention.
class foo;
  localparam int Hello_World = 1;
endclass
