`include "included-file-1.svh"

//- @MyClassIncludedFile2 defines/binding MyClassIncludedFile2
class MyClassIncludedFile2;
    //- @var5 defines/binding Var5
    static int var5;

    //- @my_fun3 defines/binding MyFun3
    function int my_fun3();
        //- @var6 ref Var6
        return var6;
    endfunction
endclass
