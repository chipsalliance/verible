`define FOO(arg) "foo``arg``bar"
