package endif_comment;
`ifdef FOOBAR
  localparam int P = 4;
`endif
endpackage
