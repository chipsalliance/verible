function foo();
endfunction
