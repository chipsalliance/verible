package does_not_match_filename_pkg;
endpackage
