module suggest_parentheses_example;
  assign foo = condition_a? condition_b? a : b : c;
endmodule
