task automatic foo;
  $psprintf("use $display\n");
endtask
