// Expected parameter type name, "Hello_World" to follow lower_snake_case naming convention and end with _t.
parameter type Hello_World = logic;
