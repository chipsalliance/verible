module posix_eof; endmodule