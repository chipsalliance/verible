// should be [0:3] or [4] according to style
logic foo [3:0];
