package endif_comment_pkg;
`ifdef FOOBAR
  parameter int P = 4;
`endif
endpackage
