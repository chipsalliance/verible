// Enum names should be lower_snake_case and end with '_t' or '_e'
typedef enum {
    Idle, Busy
} camelEnum;
