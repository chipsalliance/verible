//- @c1 defines/binding _
class c1;

    //- @var1 defines/binding _
    shortreal var1;

    //- @var2 defines/binding _
    event var2;
    
    //- @var3 defines/binding _
    chandle var3;

    //- @var4 defines/binding _
    realtime var4;

    //- @var5 defines/binding _
    real var5;

    //- @var6 defines/binding _
    int var6;

    //- @var7 defines/binding _
    logic var7;

    //- @var8 defines/binding _
    bit var8;

    //- @var9 defines/binding _
    string var9;

endclass
