// verilog_syntax: parse-as-module-body
genvar k;
for (k = 0; k < FooParam; k++) begin : gen_loop
  // code
end
