// Copyright 2020 Google LLC.
// SPDX-License-Identifier: Apache-2.0

//- @B defines/binding B
//- @A ref A
localparam B = A + 1;
