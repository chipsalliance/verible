module trailing_spaces;
endmodule 
