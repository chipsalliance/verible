module always_comb_blocking;
  always_comb
    a <= b; // [Style: combinational-logic] [always-comb-blocking]
endmodule
