// should be [3:0] according to style
logic [0:3] foo;
