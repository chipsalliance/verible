module always_comb_blocking;
  always_comb begin
    a <= b; // [Style: combinational-logic] [always-comb-blocking]
  end
endmodule
