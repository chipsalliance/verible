// verilog_syntax: parse-as-module-body
wire foo;
bar baz(x, y, z);
