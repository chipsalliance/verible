// verilog_syntax: parse-as-module-body
// Test the integration of excerpt-parsing with lint-waiving.
// This test case should trigger a line-length violation without a waiver.
assign x = f;
assign lllllllllllllllllll[1111111111] = aaaaaaaaaaa[4444444].ffffffffffffff.gggggggggggg.hhhhhhhhhhh.wwwww[555555].zzzzzzzzzz;
