//- @bad_goal ref _
module bad_goal;
endmodule
