module ILLEGALNAME; endmodule
