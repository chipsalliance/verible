module suggest_parentheses_example;
  wire foo;

  assign foo = condition_a? condition_b? a : b : c;
endmodule
