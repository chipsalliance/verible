// verilog_syntax: parse-as-module-body
generate if (foo) begin
  baz bam;
end
endgenerate
