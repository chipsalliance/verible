class foo;
  function bar;
    // The use of $test$plusargs() is not allowed.
    if ($test$plusargs("baz")) return 1;
  endfunction
endclass
